
/// This is mostly used for testing the static guarantees currently.
/// A realistic implementation would probably take four cycles.
module pipelined_mult (
    input wire clk,
    input wire reset,
    // inputs
    input wire [31:0] left,
    input wire [31:0] right,
    // The input has been committed
    output wire [31:0] out
);

logic [31:0] lt, rt, buff0, buff1, buff2, tmp_prod;

assign out = buff2;
assign tmp_prod = lt * rt;

always_ff @(posedge clk) begin
    if (reset) begin
        lt <= 0;
        rt <= 0;
        buff0 <= 0;
        buff1 <= 0;
        buff2 <= 0;
    end else begin
        lt <= left;
        rt <= right;
        buff0 <= tmp_prod;
        buff1 <= buff0;
        buff2 <= buff1;
    end
end

endmodule

module bb_pipelined_mult(
	               input wire [31:0] left,
	               input wire [31:0] right,
	               output wire [31:0] out,
	               input wire clk
	               );
`ifdef __ICARUS__
   reg [31:0] reg0;
   reg [31:0] reg1;
   reg [31:0] reg2;
   reg [31:0] reg3;
   always @( posedge clk ) begin
      reg0 <= left * right;
      reg1 <= reg0;
      reg2 <= reg1;
      reg3 <= reg2;
   end
   assign out = reg3;
`elsif VERILATOR
   reg [31:0] reg0;
   reg [31:0] reg1;
   reg [31:0] reg2;
   reg [31:0] reg3;
   always @( posedge clk ) begin
      reg0 <= left * right;
      reg1 <= reg0;
      reg2 <= reg1;
      reg3 <= reg2;
   end
   assign out = reg3;
`else
   // mul_uint32 is a black box module generated by Xilinx's IP Core generator.
   // Generation commands are in the synth.tcl file.
   mul_uint32 mul_uint32 (
                   .A(left),
                   .B(right),
                   .P(out),
                   .CLK(clk)
                   );
`endif
endmodule